// Multiplication operators between two floating-point numbers
module MultiOp (
    output [31:0] out,
    output under_overflow,
    input [31:0] para1,
    input [31:0] para2
);
// initialize variables


// mutiply fraction elements

// calculate exponent parts


//
endmodule