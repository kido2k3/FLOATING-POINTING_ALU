// the top module

module FP_ALU (
    output [31:0] out,
    output under_overflow,
    output zero,
    input [31:0] para1,
    input [31:0] para2,
    input [1:0] ALU_op
);
// initialize variables


endmodule