// Subtraction operators between two floating-point numbers
module SubOp (
    output [31:0] out,
    output under_overflow,
    input [31:0] para1,
    input [31:0] para2
);
// initialize variables


endmodule